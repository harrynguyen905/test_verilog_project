testbencc